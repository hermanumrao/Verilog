module invert(input wire i, output wire o1);
	Write code here
endmodule

module and2(input wire i0, i1, output wire o2);
	Write code here
endmodule

module or2(input wire i0, i1, output wire o3);
	Write code here
endmodule

module xor2(input wire i0, i1, output wire o4);
	Write code here
endmodule

module nand2(input wire i0, i1, output wire o5);
	wire t;
	Write code here
endmodule
