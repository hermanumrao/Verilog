module mux4 (input wire [0:3] i, input wire j1, j0, output wire o);
  wire  t0, t1;
  
Write your code here (Use only 2:1 Mux)

endmodule

